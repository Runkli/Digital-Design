library verilog;
use verilog.vl_types.all;
entity ripplecarry_vlg_vec_tst is
end ripplecarry_vlg_vec_tst;
