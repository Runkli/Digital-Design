library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity ripplecarry is
 Port (cin : in STD_LOGIC;
		 x : in STD_LOGIC_VECTOR (3 downto 0);
		 y : in STD_LOGIC_VECTOR (3 downto 0);
		 s : out STD_LOGIC_VECTOR (3 downto 0);
		 cout : out STD_LOGIC);
end ripplecarry;

architecture Structure of ripplecarry is
-- declare internal signals used to interconnect 1-bit adders:
	signal c1, c2, c3 : STD_LOGIC;
-- declare the component to be used in this architecture:
component add1bit
	 Port ( cin : in STD_LOGIC;
		 a : in STD_LOGIC;
		 b : in STD_LOGIC;
		 cout : out STD_LOGIC;
		 sum : out STD_LOGIC);
end component;

begin
-- Instantiate 1-bit adder four times and interconnect:
	stage0: add1bit port map(cin,x(0),y(0),c1,s(0));
	stage1: add1bit port map(c1,x(1),y(1),c2,s(1));
	stage2: add1bit port map(c2,x(2),y(2),c3,s(2));
	stage3: add1bit port map(c3,x(3),y(3),cout,s(3));
end Structure;
