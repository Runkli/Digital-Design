library verilog;
use verilog.vl_types.all;
entity hexdecoder_vlg_vec_tst is
end hexdecoder_vlg_vec_tst;
